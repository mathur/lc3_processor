library verilog;
use verilog.vl_types.all;
entity dcache_datapath_sv_unit is
end dcache_datapath_sv_unit;
