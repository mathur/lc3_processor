library verilog;
use verilog.vl_types.all;
entity ex_datapath_sv_unit is
end ex_datapath_sv_unit;
