library verilog;
use verilog.vl_types.all;
entity mem_io_sv_unit is
end mem_io_sv_unit;
