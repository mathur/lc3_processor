import lc3b_types::*;

module wb_datapath (
    input clk
);

endmodule : wb_datapath