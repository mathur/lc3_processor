library verilog;
use verilog.vl_types.all;
entity cache_block_sv_unit is
end cache_block_sv_unit;
