library verilog;
use verilog.vl_types.all;
entity id_datapath_sv_unit is
end id_datapath_sv_unit;
