library verilog;
use verilog.vl_types.all;
entity cpu_datapath_sv_unit is
end cpu_datapath_sv_unit;
