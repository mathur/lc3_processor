import lc3b_types::*;

module cpu_datapath
(
    input clk
);

endmodule : cpu_datapath