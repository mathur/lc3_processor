library verilog;
use verilog.vl_types.all;
entity cpu_sv_unit is
end cpu_sv_unit;
