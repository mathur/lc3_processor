library verilog;
use verilog.vl_types.all;
entity dcache_sv_unit is
end dcache_sv_unit;
