library verilog;
use verilog.vl_types.all;
entity l2_cache_sv_unit is
end l2_cache_sv_unit;
