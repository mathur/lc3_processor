library verilog;
use verilog.vl_types.all;
entity adjns_sv_unit is
end adjns_sv_unit;
