library verilog;
use verilog.vl_types.all;
entity byte_insert_sv_unit is
end byte_insert_sv_unit;
