library verilog;
use verilog.vl_types.all;
entity dcache_control_sv_unit is
end dcache_control_sv_unit;
