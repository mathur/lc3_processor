library verilog;
use verilog.vl_types.all;
entity mem_datapath_sv_unit is
end mem_datapath_sv_unit;
