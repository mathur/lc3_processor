library verilog;
use verilog.vl_types.all;
entity cache_set_sv_unit is
end cache_set_sv_unit;
