library verilog;
use verilog.vl_types.all;
entity leap_frog_sv_unit is
end leap_frog_sv_unit;
