library verilog;
use verilog.vl_types.all;
entity cache_sv_unit is
end cache_sv_unit;
