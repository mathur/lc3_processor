library verilog;
use verilog.vl_types.all;
entity if_datapath_sv_unit is
end if_datapath_sv_unit;
