library verilog;
use verilog.vl_types.all;
entity udjns_sv_unit is
end udjns_sv_unit;
