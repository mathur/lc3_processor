library verilog;
use verilog.vl_types.all;
entity udj_sv_unit is
end udj_sv_unit;
