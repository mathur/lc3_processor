library verilog;
use verilog.vl_types.all;
entity buffer_sv_unit is
end buffer_sv_unit;
