library verilog;
use verilog.vl_types.all;
entity lru_sv_unit is
end lru_sv_unit;
