library verilog;
use verilog.vl_types.all;
entity arbiter_sv_unit is
end arbiter_sv_unit;
